module rv32i_bitmap16by12(rst, clk, we, cs, addr, out);
input rst, clk, we, cs;
input [31:0] addr;
output [31:0] out;
reg [31:0] out;
reg [255:0] chr [127:0];

localparam chr_space = 7'd32;
localparam chr_excl = 7'd33;
localparam chr_dquote = 7'd34;
localparam chr_sharp = 7'd35;
localparam chr_dollar = 7'd36;
localparam chr_perc = 7'd37;
localparam chr_and = 7'd38;
localparam chr_squote = 7'd39;
localparam chr_lpar = 7'd40;
localparam chr_rpar = 7'd41;
localparam chr_star = 7'd42;
localparam chr_plus = 7'd43;
localparam chr_comma = 7'd44;
localparam chr_hyphen = 7'd45;
localparam chr_period = 7'd46;
localparam chr_fslash = 7'd47;
localparam chr_0 = 7'd48;
localparam chr_1 = 7'd49;
localparam chr_2 = 7'd50;
localparam chr_3 = 7'd51;
localparam chr_4 = 7'd52;
localparam chr_5 = 7'd53;
localparam chr_6 = 7'd54;
localparam chr_7 = 7'd55;
localparam chr_8 = 7'd56;
localparam chr_9 = 7'd57;
localparam chr_colon = 7'd58;
localparam chr_scolon = 7'd59;
localparam chr_lthan = 7'd60;
localparam chr_equal = 7'd61;
localparam chr_gthan = 7'd62;
localparam chr_ques = 7'd63;
localparam chr_at = 7'd64;
localparam chr_A = 7'd65;
localparam chr_B = 7'd66;
localparam chr_C = 7'd67;
localparam chr_D = 7'd68;
localparam chr_E = 7'd69;
localparam chr_F = 7'd70;
localparam chr_G = 7'd71;
localparam chr_H = 7'd72;
localparam chr_I = 7'd73;
localparam chr_J = 7'd74;
localparam chr_K = 7'd75;
localparam chr_L = 7'd76;
localparam chr_M = 7'd77;
localparam chr_N = 7'd78;
localparam chr_O = 7'd79;
localparam chr_P = 7'd80;
localparam chr_Q = 7'd81;
localparam chr_R = 7'd82;
localparam chr_S = 7'd83;
localparam chr_T = 7'd84;
localparam chr_U = 7'd85;
localparam chr_V = 7'd86;
localparam chr_W = 7'd87;
localparam chr_X = 7'd88;
localparam chr_Y = 7'd89;
localparam chr_Z = 7'd90;
localparam chr_lbrack = 7'd91;
localparam chr_bslash = 7'd92;
localparam chr_rbrack = 7'd93;
localparam chr_exp = 7'd94;
localparam chr_uscore = 7'd95;
localparam chr_apo = 7'd96;
localparam chr_a = 7'd97;
localparam chr_b = 7'd98;
localparam chr_c = 7'd99;
localparam chr_d = 7'd100;
localparam chr_e = 7'd101;
localparam chr_f = 7'd102;
localparam chr_g = 7'd103;
localparam chr_h = 7'd104;
localparam chr_i = 7'd105;
localparam chr_j = 7'd106;
localparam chr_k = 7'd107;
localparam chr_l = 7'd108;
localparam chr_m = 7'd109;
localparam chr_n = 7'd110;
localparam chr_o = 7'd111;
localparam chr_p = 7'd112;
localparam chr_q = 7'd113;
localparam chr_r = 7'd114;
localparam chr_s = 7'd115;
localparam chr_t = 7'd116;
localparam chr_u = 7'd117;
localparam chr_v = 7'd118;
localparam chr_w = 7'd119;
localparam chr_x = 7'd120;
localparam chr_y = 7'd121;
localparam chr_z = 7'd122;
localparam chr_lbrace = 7'd123;
localparam chr_or = 7'd124;
localparam chr_rbrace = 7'd125;
localparam chr_wave = 7'd126;
localparam chr_del = 7'd127;

always @(posedge rst, posedge clk)
begin
	if(rst)
	begin
		chr[chr_space] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
		chr[chr_excl] <= 256'h00000000000000000000000000000000000000007FCC00000000000000000000;
		chr[chr_dquote] <= 256'h0000000000000000000000000000000078000000000078000000000000000000;
		chr[chr_sharp] <= 256'h000000000000000000000000024002401FF8024002401FF80240024000000000;
		chr[chr_dollar] <= 256'h00000000000000000000000010602090210821087FFC210812080C1000000000;
		chr[chr_perc] <= 256'h000000000000000000000000000030180C24031800C01830240C180000000000;
		chr[chr_and] <= 256'h00000000000000000000000000403C44424842B0410842043D0800F000000000;
		chr[chr_squote] <= 256'h0000000000000000000000000000000000000000780000000000000000000000;
		chr[chr_lpar] <= 256'h000000000000000000000000000000000000600C183007C00000000000000000;
		chr[chr_rpar] <= 256'h0000000000000000000000000000000007C01830600C00000000000000000000;
		chr[chr_star] <= 256'h00000000000000000000000000000000008006B001C001C006B0008000000000;
		chr[chr_plus] <= 256'h000000000000000000000000000000800080008007F000800080008000000000;
		chr[chr_comma] <= 256'h0000000000000000000000000000000000000030000C00000000000000000000;
		chr[chr_hyphen] <= 256'h0000000000000000000000000000010001000100010001000100000000000000;
		chr[chr_period] <= 256'h0000000000000000000000000000000000000000000C000C0000000000000000;
		chr[chr_fslash] <= 256'h000000000000000000000000000030000C00030000C00030000C000000000000;
		chr[chr_0] <= 256'h0000000000000000000000001FF02008400441844184400420081FF000000000;
		chr[chr_1] <= 256'h00000000000000000000000000000000000400047FFC30041004000000000000;
		chr[chr_2] <= 256'h0000000000000000000000001C04220441044084404440242014180C00000000;
		chr[chr_3] <= 256'h00000000000000000000000000F03D0842044204420440042008101000000000;
		chr[chr_4] <= 256'h00000000000000000000000000807FFC20801080088004800280018000000000;
		chr[chr_5] <= 256'h00000000000000000000000041F04208440444044404440442047E0400000000;
		chr[chr_6] <= 256'h00000000000000000000000010F02108420442044204420423081FF000000000;
		chr[chr_7] <= 256'h00000000000000000000000070004C00430040C04030400C4000400000000000;
		chr[chr_8] <= 256'h00000000000000000000000000F03D0842044204420442043D0800F000000000;
		chr[chr_9] <= 256'h0000000000000000000000001FF02108408440844084408421081E1000000000;
		chr[chr_colon] <= 256'h0000000000000000000000000000000000000660066000000000000000000000;
		chr[chr_scolon] <= 256'h0000000000000000000000000000000000000660061800000000000000000000;
		chr[chr_lthan] <= 256'h0000000000000000000000000810081004200420024002400180018000000000;
		chr[chr_equal] <= 256'h0000000000000000000000000240024002400240024002400240000000000000;
		chr[chr_gthan] <= 256'h0000000000000000000001800180024002400420042008100810000000000000;
		chr[chr_ques] <= 256'h0000000000000000000000001E0021004080404C404C40002000180000000000;
		chr[chr_at] <= 256'h0000000000000000000000001F9020484FE44824482447C420081FF000000000;
		chr[chr_A] <= 256'h0000000000000000000000003FFC4080408040804080408040803FFC00000000;
		chr[chr_B] <= 256'h00000000000000000000000018F02508420442044204420442047FFC00000000;
		chr[chr_C] <= 256'h00000000000000000000000040044004400440044004400420081FF000000000;
		chr[chr_D] <= 256'h0000000000000000000000001FF02008400440044004400440047FFC00000000;
		chr[chr_E] <= 256'h00000000000000000000000040044004400442044204420442047FFC00000000;
		chr[chr_F] <= 256'h00000000000000000000000040004000400042004200420042007FFC00000000;
		chr[chr_G] <= 256'h00000000000000000000000021F04108410441044004400420081FF000000000;
		chr[chr_H] <= 256'h0000000000000000000000007FFC0100010001000100010001007FFC00000000;
		chr[chr_I] <= 256'h00000000000000000000000000000000400440047FFC40044004000000000000;
		chr[chr_J] <= 256'h0000000000000000000000007FF0400840044004400440044004400400000000;
		chr[chr_K] <= 256'h00000000000000000000000040042008101008200440028001007FFC00000000;
		chr[chr_L] <= 256'h00000000000000000000000000040004000400040004000400047FFC00000000;
		chr[chr_M] <= 256'h0000000000000000000000007FFC30000C00020002000C0030007FFC00000000;
		chr[chr_N] <= 256'h0000000000000000000000007FFC001C006001800600180060007FFC00000000;
		chr[chr_O] <= 256'h0000000000000000000000001FF02008400440044004400420081FF000000000;
		chr[chr_P] <= 256'h0000000000000000000000001E002100408040804080408040807FFC00000000;
		chr[chr_Q] <= 256'h0000000000000000000000001FEC2018403C40644004400420081FF000000000;
		chr[chr_R] <= 256'h0000000000000000000000001E042108409040A040C0408040807FFC00000000;
		chr[chr_S] <= 256'h00000000000000000000000000702088410441044104410422081C0000000000;
		chr[chr_T] <= 256'h00000000000000000000000040004000400040007FFC40004000400000000000;
		chr[chr_U] <= 256'h0000000000000000000000007FF00008000400040004000400087FF000000000;
		chr[chr_V] <= 256'h0000000000000000000000007800070000E0001C001C00E00700780000000000;
		chr[chr_W] <= 256'h0000000000000000000000007F80007C001807E007E00018007C7F8000000000;
		chr[chr_X] <= 256'h000000000000000000000000600C183006C00100010006C01830600C00000000;
		chr[chr_Y] <= 256'h00000000000000000000000060001800060001FC01FC06001800600000000000;
		chr[chr_Z] <= 256'h0000000000000000000000006004580446044104410440C44034400C00000000;
		chr[chr_lbrack] <= 256'h000000000000000000000000000000004004400440047FFC0000000000000000;
		chr[chr_bslash] <= 256'h0000000000000000000000000000000C003000C003000C003000000000000000;
		chr[chr_rbrack] <= 256'h000000000000000000000000000000007FFC4004400440040000000000000000;
		chr[chr_exp] <= 256'h0000000000000000000000000800100020004000400020001000080000000000;
		chr[chr_uscore] <= 256'h0000000000000000000000000004000400040004000400040004000400000000;
		chr[chr_apo] <= 256'h0000000000000000000000000000000000001800600000000000000000000000;
		chr[chr_a] <= 256'h00000000000000000000000003FC01080204020402040204010800F000000000;
		chr[chr_b] <= 256'h00000000000000000000000000F00108020402040204020402047FFC00000000;
		chr[chr_c] <= 256'h000000000000000000000000010802040204020402040204010800F000000000;
		chr[chr_d] <= 256'h0000000000000000000000007FFC02040204020402040204010800F000000000;
		chr[chr_e] <= 256'h00000000000000000000000001C802440244024402440244014800F000000000;
		chr[chr_f] <= 256'h0000000000000000000000000000400040004000400020801FFC008000000000;
		chr[chr_g] <= 256'h00000000000000000000000003F0044808440844084408440484030800000000;
		chr[chr_h] <= 256'h000000000000000000000000007C0080010001000100010001007FFC00000000;
		chr[chr_i] <= 256'h0000000000000000000000000000000000000000037C00000000000000000000;
		chr[chr_j] <= 256'h00000000000000000000000000000000000006F0000800040000000000000000;
		chr[chr_k] <= 256'h00000000000000000000000001040104008800880050005000207FFC00000000;
		chr[chr_l] <= 256'h000000000000000000000000000000000004000400047FF80000000000000000;
		chr[chr_m] <= 256'h00000000000000000000000001FC0200010000C000C00100020001FC00000000;
		chr[chr_n] <= 256'h00000000000000000000000001FC02000200020002000200020001FC00000000;
		chr[chr_o] <= 256'h00000000000000000000000000F001080204020402040204010800F000000000;
		chr[chr_p] <= 256'h00000000000000000000000003000480084008400840084008400FFC00000000;
		chr[chr_q] <= 256'h0000000000000000000000000FFC084008400840084008400480030000000000;
		chr[chr_r] <= 256'h00000000000000000000000000000200020002000100010003FC000000000000;
		chr[chr_s] <= 256'h0000000000000000000000000110022804440444044404440288011000000000;
		chr[chr_t] <= 256'h00000000000000000000000000000000080008007FFC08000800000000000000;
		chr[chr_u] <= 256'h00000000000000000000000003FC00080004000400040004000803F000000000;
		chr[chr_v] <= 256'h000000000000000000000000030000C00030000C000C003000C0030000000000;
		chr[chr_w] <= 256'h00000000000000000000000003C0003C0010007000700010003C03C000000000;
		chr[chr_x] <= 256'h0000000000000000000000000204010800900060006000900108020400000000;
		chr[chr_y] <= 256'h0000000000000000000000000200010000800078004400840104020000000000;
		chr[chr_z] <= 256'h0000000000000000000000000304028402440244022402240214020C00000000;
		chr[chr_lbrace] <= 256'h00000000000000000000000000004004400420081EF001000100000000000000;
		chr[chr_or] <= 256'h00000000000000000000000000000000000000007FFC00000000000000000000;
		chr[chr_rbrace] <= 256'h0000000000000000000000000000010001001EF0200840044004000000000000;
		chr[chr_wave] <= 256'h0000000000000000000000000180004000400080010002000200018000000000;
		chr[chr_del] <= 256'h00000000000000000000010001000100010001000100010007c0038001000000;
		out <= 32'bz;
	end
	else
	begin
		if((cs==1)&&(we==0)&&(addr[31:12]>=20'hE0001)&&(addr[31:12]<=20'hE000F)) //
		begin
			out[31:16] <= 0;
			case(addr[4:1])
			4'b0000: out[15:0] <= chr[addr[11:5]][0*16+15:0*16]; //column 0
			4'b0001: out[15:0] <= chr[addr[11:5]][1*16+15:1*16]; //column 1
		   4'b0010: out[15:0] <= chr[addr[11:5]][2*16+15:2*16]; 
			4'b0011: out[15:0] <= chr[addr[11:5]][3*16+15:3*16];
			4'b0100: out[15:0] <= chr[addr[11:5]][4*16+15:4*16];
			4'b0101: out[15:0] <= chr[addr[11:5]][5*16+15:5*16];
			4'b0110: out[15:0] <= chr[addr[11:5]][6*16+15:6*16];
			4'b0111: out[15:0] <= chr[addr[11:5]][7*16+15:7*16];
			4'b1000: out[15:0] <= chr[addr[11:5]][8*16+15:8*16];
			4'b1001: out[15:0] <= chr[addr[11:5]][9*16+15:9*16];
		   4'b1010: out[15:0] <= chr[addr[11:5]][10*16+15:10*16];
			4'b1011: out[15:0] <= chr[addr[11:5]][11*16+15:11*16]; //column 11
			4'b1100: out[15:0] <= chr[addr[11:5]][12*16+15:12*16]; //unused
			4'b1101: out[15:0] <= chr[addr[11:5]][13*16+15:13*16]; //unused
			4'b1110: out[15:0] <= chr[addr[11:5]][14*16+15:14*16]; //unused
			4'b1111: out[15:0] <= chr[addr[11:5]][15*16+15:15*16]; //unused
			endcase
		end
		else out <= 32'bz;
	end
end

endmodule
